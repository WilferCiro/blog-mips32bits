// Wilfer Daniel Ciro Maya - 2023

module flash(dir, opCode);
	// parameters definitions
	parameter BUS_SIZE = 32;
	parameter DIR_SIZE = 32;
	parameter OPC_SIZE = BUS_SIZE;
	
	parameter MEM_SIZE = 255;
	
	// inputs declarations
	input [DIR_SIZE - 1 : 0] dir;
	
	// outputs declarations
	output [OPC_SIZE - 1 : 0] opCode;
	
	// firmware, change for the correct firmware to exec
	reg [OPC_SIZE - 1 : 0] ROM [0 : MEM_SIZE];
	initial
	begin
		//$readmemb("/home/ciro/Documents/Universidad/Semestre9/DDA/ROMMicro.mem", ROM);
		
		ROM[0] = 32'b001111_00000_00001_00000_00000000001; // LUI reg1 = 1 -> para asignar a la salida
		// Assign ports positions
		ROM[1] = 32'b001111_00000_00010_00000_00000000010; // LUI reg2 = 2
		ROM[2] = 32'b001111_00000_00011_00000_00000000011; // LUI reg3 = 3
		ROM[3] = 32'b001111_00000_00100_00000_00000000100; // LUI reg4 = 4
		ROM[4] = 32'b001111_00000_00101_00000_00000000101; // LUI reg5 = 5
		ROM[5] = 32'b001111_00000_00110_00000_00000000110; // LUI reg6 = 6
		ROM[6] = 32'b001111_00000_00111_00000_00000000111; // LUI reg7 = 7
		
		
		ROM[7] = 32'b001111_00000_01000_00000_00000001000; // LUI reg8 = 8 -> pin entrada 8
		ROM[8] = 32'b001111_00000_01001_00000_00000001001; // LUI reg9 = 9 -> pin entrada 8
		ROM[9] = 32'b001111_00000_10001_00000_00000000000; // LUI reg17 = 0 -> para sumar de 0 - 9
		
		ROM[10] = 32'b001111_00000_11010_00000_00000000000; // LUI reg26 = 0 -> para sumar de 0 - 9
				
		/* DELAY TIME */
		ROM[11] = 32'b001111_00000_01011_01111_11111111111; // LUI reg11 = max -> para delay
		
		ROM[12] = 32'b001111_00000_10101_00000_00000000000; // LUI reg21 = 0 -> para delay
		ROM[13] = 32'b001111_00000_10110_00000_00001111111; // LUI reg22 = 21 -> para delay		
		ROM[14] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[15] = 32'b000000_00000_00000_00000_00000000000; // NOP		
		ROM[16] = 32'b001000_10101_10101_00000_00000000001; // reg21 ++	
		ROM[17] = 32'b001000_01011_01011_01111_11111111111; // Reg11 += Reg11
		ROM[18] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[19] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[20] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[21] = 32'b000100_10101_10110_0000000000000011; // BEQ reg21 == reg22 (2) -> Ir a encender
		ROM[22] = 32'b000010_11111_11111_1111111111111001; // Jump (-7)	
		ROM[23] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
	
		/* IDLE */
		ROM[24] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[25] = 32'b000000_00000_00000_00000_00000000000; // NOP		
		ROM[26] = 32'b100011_01000_10000_00000_00000000000; // Reg16 = read_pin_8 (reg2)
		ROM[27] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[28] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[29] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[30] = 32'b000100_00001_10000_0000000000000100; // BEQ reg1 == reg16 (3) -> ir a aumentar
		ROM[31] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[32] = 32'b000010_11111_11111_1111111111111001; // Jump (-7)
		ROM[33] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		/* DELAY */
		ROM[34] = 32'b001111_00000_01010_00000_00000000000; // LUI reg10 = 0 -> para delay		
		
		ROM[35] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[36] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[37] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		ROM[38] = 32'b001000_01010_01010_00000_00000000001; // Reg10 ++
		
		ROM[39] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[40] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[41] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[42] = 32'b000100_01011_01010_0000000000000011; // BEQ reg10 == reg11 (2) -> Ir a encender
		ROM[43] = 32'b000010_11111_11111_1111111111111001; // Jump (-7)	
		ROM[44] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		/*	Aumentar y Encender */
		ROM[45] = 32'b001000_10001_10001_00000_00000000001; // Reg17 ++		
		ROM[46] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[47] = 32'b000000_00000_00000_00000_00000000000; // NOP
		ROM[48] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// if 0
		ROM[49] = 32'b000100_00000_10001_0000000000010100; // BEQ reg17 == reg0 (20) / enciende 0
		ROM[50] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// if 1
		ROM[51] = 32'b000100_00001_10001_0000000000011011; // BEQ reg17 == reg1 (27) / enciende 1
		ROM[52] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// if 2
		ROM[53] = 32'b000100_00010_10001_0000000000100010; // BEQ reg17 == reg2 (34) / enciende 2
		ROM[54] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// if 3
		ROM[55] = 32'b000100_00011_10001_0000000000101001; // BEQ reg17 == reg3 (41) / enciende 3
		ROM[56] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// if 4
		ROM[57] = 32'b000100_00100_10001_0000000000110000; // BEQ reg17 == reg4 (48) / enciende 3
		ROM[58] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// if 5
		ROM[59] = 32'b000100_00101_10001_0000000000110111; // BEQ reg17 == reg5 (55) / enciende 3
		ROM[60] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// if 6
		ROM[61] = 32'b000100_00110_10001_0000000000111110; // BEQ reg17 == reg6 (62) / enciende 3
		ROM[62] = 32'b000000_00000_00000_00000_00000000000; // NOP
	
		// if 7
		ROM[63] = 32'b000100_00111_10001_0000000001000101; // BEQ reg17 == reg7 (69) / enciende 3
		ROM[64] = 32'b000000_00000_00000_00000_00000000000; // NOP
	
		// if 8
		ROM[65] = 32'b000100_01000_10001_0000000001001100; // BEQ reg17 == reg8 (76) / enciende 3
		ROM[66] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// if 9
		ROM[67] = 32'b000100_01001_10001_0000000001010011; // BEQ reg17 == reg9 (83) / enciende 3
		ROM[68] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
				
		/* Encender */
		// el 0
		ROM[69] = 32'b101011_00000_00001_00000_00000000000; // port0 = reg1
		ROM[70] = 32'b101011_00001_00001_00000_00000000000; // port1 = reg1
		ROM[71] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[72] = 32'b101011_00011_00001_00000_00000000000; // port3 = reg1
		ROM[73] = 32'b101011_00100_00001_00000_00000000000; // port4 = reg1
		ROM[74] = 32'b101011_00101_00001_00000_00000000000; // port5 = reg1
		ROM[75] = 32'b101011_00110_00000_00000_00000000000; // port6 = reg0
		
		ROM[76] = 32'b000010_11111_11111_1111111111001100; // Jump (-52)
			
		ROM[77] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// el 1
		ROM[78] = 32'b101011_00000_00000_00000_00000000000; // port0 = reg0
		ROM[79] = 32'b101011_00001_00001_00000_00000000000; // port1 = reg0
		ROM[80] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[81] = 32'b101011_00011_00000_00000_00000000000; // port3 = reg1
		ROM[82] = 32'b101011_00100_00000_00000_00000000000; // port4 = reg1
		ROM[83] = 32'b101011_00101_00000_00000_00000000000; // port5 = reg1
		ROM[84] = 32'b101011_00110_00000_00000_00000000000; // port6 = reg1		
		ROM[85] = 32'b000010_11111_11111_1111111111000011; // Jump (-61)			
		ROM[86] = 32'b000000_00000_00000_00000_00000000000; // NOP
	
		// el 2
		ROM[87] = 32'b101011_00000_00001_00000_00000000000; // port7 = reg0
		ROM[88] = 32'b101011_00001_00001_00000_00000000000; // port1 = reg0
		ROM[89] = 32'b101011_00010_00000_00000_00000000000; // port2 = reg1
		ROM[90] = 32'b101011_00011_00001_00000_00000000000; // port3 = reg1
		ROM[91] = 32'b101011_00100_00001_00000_00000000000; // port4 = reg1
		ROM[92] = 32'b101011_00101_00000_00000_00000000000; // port5 = reg1
		ROM[93] = 32'b101011_00110_00001_00000_00000000000; // port6 = reg1
		
		ROM[94] = 32'b000010_11111_11111_1111111110111010; // Jump (-70)
			
		ROM[95] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// el 3
		ROM[96] = 32'b101011_00000_00001_00000_00000000000; // port7 = reg0
		ROM[97] = 32'b101011_00001_00001_00000_00000000000; // port1 = reg0
		ROM[98] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[99] = 32'b101011_00011_00001_00000_00000000000; // port3 = reg1
		ROM[100] = 32'b101011_00100_00000_00000_00000000000; // port4 = reg1
		ROM[101] = 32'b101011_00101_00000_00000_00000000000; // port5 = reg1
		ROM[102] = 32'b101011_00110_00001_00000_00000000000; // port6 = reg1		
		ROM[103] = 32'b000010_11111_11111_1111111110110001; // Jump (-79)			
		ROM[104] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// el 4
		ROM[105] = 32'b101011_00000_00000_00000_00000000000; // port7 = reg0
		ROM[106] = 32'b101011_00001_00001_00000_00000000000; // port1 = reg0
		ROM[107] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[108] = 32'b101011_00011_00000_00000_00000000000; // port3 = reg1
		ROM[109] = 32'b101011_00100_00000_00000_00000000000; // port4 = reg1
		ROM[110] = 32'b101011_00101_00001_00000_00000000000; // port5 = reg1
		ROM[111] = 32'b101011_00110_00001_00000_00000000000; // port6 = reg1
		ROM[112] = 32'b000010_11111_11111_1111111110101000; // Jump (-88)			
		ROM[113] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// el 5
		ROM[114] = 32'b101011_00000_00001_00000_00000000000; // port7 = reg0
		ROM[115] = 32'b101011_00001_00000_00000_00000000000; // port1 = reg0
		ROM[116] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[117] = 32'b101011_00011_00001_00000_00000000000; // port3 = reg1
		ROM[118] = 32'b101011_00100_00000_00000_00000000000; // port4 = reg1
		ROM[119] = 32'b101011_00101_00001_00000_00000000000; // port5 = reg1
		ROM[120] = 32'b101011_00110_00001_00000_00000000000; // port6 = reg1		
		ROM[121] = 32'b000010_11111_11111_1111111110011111; // Jump (-97)			
		ROM[122] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// el 6
		ROM[123] = 32'b101011_00000_00001_00000_00000000000; // port7 = reg0
		ROM[124] = 32'b101011_00001_00000_00000_00000000000; // port1 = reg0
		ROM[125] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[126] = 32'b101011_00011_00001_00000_00000000000; // port3 = reg1
		ROM[127] = 32'b101011_00100_00001_00000_00000000000; // port4 = reg1
		ROM[128] = 32'b101011_00101_00001_00000_00000000000; // port5 = reg1
		ROM[129] = 32'b101011_00110_00001_00000_00000000000; // port6 = reg1		
		ROM[130] = 32'b000010_11111_11111_1111111110010110; // Jump (-106)			
		ROM[131] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// el 7
		ROM[132] = 32'b101011_00000_00001_00000_00000000000; // port7 = reg0
		ROM[133] = 32'b101011_00001_00001_00000_00000000000; // port1 = reg0
		ROM[134] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[135] = 32'b101011_00011_00000_00000_00000000000; // port3 = reg1
		ROM[136] = 32'b101011_00100_00000_00000_00000000000; // port4 = reg1
		ROM[137] = 32'b101011_00101_00000_00000_00000000000; // port5 = reg1
		ROM[138] = 32'b101011_00110_00000_00000_00000000000; // port6 = reg1		
		ROM[139] = 32'b000010_11111_11111_1111111110001101; // Jump (-115)			
		ROM[140] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// el 8
		ROM[141] = 32'b101011_00000_00001_00000_00000000000; // port7 = reg0
		ROM[142] = 32'b101011_00001_00001_00000_00000000000; // port1 = reg0
		ROM[143] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[144] = 32'b101011_00011_00001_00000_00000000000; // port3 = reg1
		ROM[145] = 32'b101011_00100_00001_00000_00000000000; // port4 = reg1
		ROM[146] = 32'b101011_00101_00001_00000_00000000000; // port5 = reg1
		ROM[147] = 32'b101011_00110_00001_00000_00000000000; // port6 = reg1		
		ROM[148] = 32'b000010_11111_11111_1111111110000100; // Jump (-124)			
		ROM[149] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		// el 9
		ROM[150] = 32'b101011_00000_00001_00000_00000000000; // port7 = reg0
		ROM[151] = 32'b101011_00001_00001_00000_00000000000; // port1 = reg0
		ROM[152] = 32'b101011_00010_00001_00000_00000000000; // port2 = reg1
		ROM[153] = 32'b101011_00011_00001_00000_00000000000; // port3 = reg1
		ROM[154] = 32'b101011_00100_00000_00000_00000000000; // port4 = reg1
		ROM[155] = 32'b101011_00101_00001_00000_00000000000; // port5 = reg1
		ROM[156] = 32'b101011_00110_00001_00000_00000000000; // port6 = reg1		
		ROM[157] = 32'b001111_00000_10001_00000_00000000000; // LUI reg17 = 0 -> para sumar de 0 - 9
					
		ROM[158] = 32'b001000_11010_11010_00000_00000000001; // Reg26 ++	
		ROM[159] = 32'b000000_00000_00000_00000_00000000000; // NOP			
		ROM[160] = 32'b000000_00000_00000_00000_00000000000; // NOP			
		ROM[161] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
		ROM[162] = 32'b101011_00111_11010_00000_00000000000; // port7 = reg26
		ROM[163] = 32'b000010_11111_11111_1111111101110101; // Jump (-135)			
		ROM[164] = 32'b000000_00000_00000_00000_00000000000; // NOP
		
	end
	/*
	integer i;
	initial begin
		for (i = 0; i <= MEM_SIZE; i = i + 1)
			ROM[i] = 32'b0;
		ROM[0] = 32'b101011_01010_000000000000001000000;
		ROM[1] = 32'b100011_01010_000000000000000010000;
		ROM[2] = 32'b101011_01010_000000000000000000100;
		ROM[3] = 32'b100010_01010_000000000000000000010;
		ROM[4] = 32'b101011_01010_000000000000001000000;
	end
	*/
	// Data flow	
	assign opCode = ROM[dir];
endmodule 
